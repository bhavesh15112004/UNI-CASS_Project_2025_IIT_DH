** sch_path: /home/designer/shared/uni_cass/final_design/Differential_ended_Design.sch
**.subckt Differential_ended_Design
V2 VDD GND 1.6
V3 v2 GND dc 0.8 ac 1
V4 v1 GND dc 0.8 ac 0
XM7 VOP nbias GND GND sg13_hv_nmos w=4u l=2u ng=1 m=1
XM8 VOP v2 tail tail sg13_hv_pmos w=9u l=1u ng=1 m=1
XM9 VOM nbias GND GND sg13_hv_nmos w=4u l=2u ng=1 m=1
XM10 VOM v1 tail tail sg13_hv_pmos w=9u l=1u ng=1 m=1
XM11 tail pbias VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=4
XM12 pbias pbias VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=1
I1 pbias GND 1u
C2 VOM GND 1p m=1
C3 VOP GND 1p m=1
XM6 net1 net1 GND GND sg13_hv_nmos w=1u l=0.5u ng=1 m=1
XM13 net1 VOP tail_cmfb tail_cmfb sg13_hv_pmos w=2.25u l=0.5u ng=1 m=1
XM14 nbias net1 GND GND sg13_hv_nmos w=1u l=0.5u ng=1 m=1
XM15 nbias VCM_REF tail_cmfb tail_cmfb sg13_hv_pmos w=4.5u l=0.5u ng=1 m=1
XM16 tail_cmfb pbias VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=4
XM17 net1 VOM tail_cmfb tail_cmfb sg13_hv_pmos w=2.25u l=0.5u ng=1 m=1
V1 VCM_REF GND dc 0.6 ac 0
C5 nbias GND 1p m=1
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ






*.ac dec 10 100 10e8
*.save all
.op



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
